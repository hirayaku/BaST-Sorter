import Vector::*;
import GetPut::*;

// a vector of Put interfaces
typedef Vector#(m, Put#(Vector#(n, itype))) Puts#(numeric type m, numeric type n, type itype);

